library verilog;
use verilog.vl_types.all;
entity altera_lnsim_functions is
end altera_lnsim_functions;
