library verilog;
use verilog.vl_types.all;
entity ama_preadder_function is
    generic(
        preadder_mode   : string  := "SIMPLE";
        width_in_a      : integer := 1;
        width_in_b      : integer := 1;
        width_in_c      : integer := 1;
        width_in_coef   : integer := 1;
        width_result_a  : integer := 1;
        width_result_b  : integer := 1;
        preadder_direction_0: string  := "ADD";
        preadder_direction_1: string  := "ADD";
        preadder_direction_2: string  := "ADD";
        preadder_direction_3: string  := "ADD";
        representation_preadder_adder: string  := "UNSIGNED";
        width_in_a_msb  : vl_notype;
        width_in_b_msb  : vl_notype;
        width_in_c_msb  : vl_notype;
        width_in_coef_msb: vl_notype;
        width_result_a_msb: vl_notype;
        width_result_b_msb: vl_notype;
        width_preadder_adder_input: vl_notype;
        width_preadder_adder_input_msb: vl_notype;
        width_preadder_adder_result: vl_notype;
        width_preadder_adder_result_msb: vl_notype;
        width_preadder_adder_input_wire: vl_notype;
        width_preadder_adder_input_wire_msb: vl_notype;
        width_in_a_ext  : vl_notype;
        width_in_b_ext  : vl_notype;
        width_output_preadder: vl_notype;
        width_output_preadder_msb: vl_notype;
        width_output_coef: vl_notype;
        width_output_coef_msb: vl_notype;
        width_output_datab: vl_notype;
        width_output_datab_msb: vl_notype;
        width_output_datac: vl_notype;
        width_output_datac_msb: vl_notype
    );
    port(
        dataa_in_0      : in     vl_logic_vector;
        dataa_in_1      : in     vl_logic_vector;
        dataa_in_2      : in     vl_logic_vector;
        dataa_in_3      : in     vl_logic_vector;
        datab_in_0      : in     vl_logic_vector;
        datab_in_1      : in     vl_logic_vector;
        datab_in_2      : in     vl_logic_vector;
        datab_in_3      : in     vl_logic_vector;
        datac_in_0      : in     vl_logic_vector;
        datac_in_1      : in     vl_logic_vector;
        datac_in_2      : in     vl_logic_vector;
        datac_in_3      : in     vl_logic_vector;
        coef0           : in     vl_logic_vector;
        coef1           : in     vl_logic_vector;
        coef2           : in     vl_logic_vector;
        coef3           : in     vl_logic_vector;
        result_a0       : out    vl_logic_vector;
        result_a1       : out    vl_logic_vector;
        result_a2       : out    vl_logic_vector;
        result_a3       : out    vl_logic_vector;
        result_b0       : out    vl_logic_vector;
        result_b1       : out    vl_logic_vector;
        result_b2       : out    vl_logic_vector;
        result_b3       : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of preadder_mode : constant is 1;
    attribute mti_svvh_generic_type of width_in_a : constant is 1;
    attribute mti_svvh_generic_type of width_in_b : constant is 1;
    attribute mti_svvh_generic_type of width_in_c : constant is 1;
    attribute mti_svvh_generic_type of width_in_coef : constant is 1;
    attribute mti_svvh_generic_type of width_result_a : constant is 1;
    attribute mti_svvh_generic_type of width_result_b : constant is 1;
    attribute mti_svvh_generic_type of preadder_direction_0 : constant is 1;
    attribute mti_svvh_generic_type of preadder_direction_1 : constant is 1;
    attribute mti_svvh_generic_type of preadder_direction_2 : constant is 1;
    attribute mti_svvh_generic_type of preadder_direction_3 : constant is 1;
    attribute mti_svvh_generic_type of representation_preadder_adder : constant is 1;
    attribute mti_svvh_generic_type of width_in_a_msb : constant is 3;
    attribute mti_svvh_generic_type of width_in_b_msb : constant is 3;
    attribute mti_svvh_generic_type of width_in_c_msb : constant is 3;
    attribute mti_svvh_generic_type of width_in_coef_msb : constant is 3;
    attribute mti_svvh_generic_type of width_result_a_msb : constant is 3;
    attribute mti_svvh_generic_type of width_result_b_msb : constant is 3;
    attribute mti_svvh_generic_type of width_preadder_adder_input : constant is 3;
    attribute mti_svvh_generic_type of width_preadder_adder_input_msb : constant is 3;
    attribute mti_svvh_generic_type of width_preadder_adder_result : constant is 3;
    attribute mti_svvh_generic_type of width_preadder_adder_result_msb : constant is 3;
    attribute mti_svvh_generic_type of width_preadder_adder_input_wire : constant is 3;
    attribute mti_svvh_generic_type of width_preadder_adder_input_wire_msb : constant is 3;
    attribute mti_svvh_generic_type of width_in_a_ext : constant is 3;
    attribute mti_svvh_generic_type of width_in_b_ext : constant is 3;
    attribute mti_svvh_generic_type of width_output_preadder : constant is 3;
    attribute mti_svvh_generic_type of width_output_preadder_msb : constant is 3;
    attribute mti_svvh_generic_type of width_output_coef : constant is 3;
    attribute mti_svvh_generic_type of width_output_coef_msb : constant is 3;
    attribute mti_svvh_generic_type of width_output_datab : constant is 3;
    attribute mti_svvh_generic_type of width_output_datab_msb : constant is 3;
    attribute mti_svvh_generic_type of width_output_datac : constant is 3;
    attribute mti_svvh_generic_type of width_output_datac_msb : constant is 3;
end ama_preadder_function;
