library verilog;
use verilog.vl_types.all;
entity altera_generic_pll_functions is
end altera_generic_pll_functions;
