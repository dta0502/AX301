library verilog;
use verilog.vl_types.all;
entity lut_input is
    port(
        \in\            : in     vl_logic;
        \out\           : out    vl_logic
    );
end lut_input;
