library verilog;
use verilog.vl_types.all;
entity ama_data_split_reg_ext_function is
    generic(
        width_data_in   : integer := 1;
        width_data_out  : vl_notype;
        register_clock_0: string  := "UNREGISTERED";
        register_aclr_0 : string  := "UNUSED";
        register_clock_1: string  := "UNREGISTERED";
        register_aclr_1 : string  := "UNUSED";
        register_clock_2: string  := "UNREGISTERED";
        register_aclr_2 : string  := "UNUSED";
        register_clock_3: string  := "UNREGISTERED";
        register_aclr_3 : string  := "UNUSED";
        number_of_multipliers: integer := 1;
        port_sign       : string  := "PORT_CONNECTIVITY";
        width_data_in_msb: vl_notype;
        width_data_in_total_msb: vl_notype;
        width_data_out_msb: vl_notype;
        width_data_in_0_msb: vl_notype;
        width_data_in_0_lsb: integer := 0;
        width_data_in_1_msb: vl_notype;
        width_data_in_1_lsb: vl_notype;
        width_data_in_2_msb: vl_notype;
        width_data_in_2_lsb: vl_notype;
        width_data_in_3_msb: vl_notype;
        width_data_in_3_lsb: vl_notype
    );
    port(
        clock           : in     vl_logic_vector(3 downto 0);
        aclr            : in     vl_logic_vector(3 downto 0);
        ena             : in     vl_logic_vector(3 downto 0);
        sign            : in     vl_logic;
        data_in         : in     vl_logic_vector;
        data_out_0      : out    vl_logic_vector;
        data_out_1      : out    vl_logic_vector;
        data_out_2      : out    vl_logic_vector;
        data_out_3      : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of width_data_in : constant is 1;
    attribute mti_svvh_generic_type of width_data_out : constant is 3;
    attribute mti_svvh_generic_type of register_clock_0 : constant is 1;
    attribute mti_svvh_generic_type of register_aclr_0 : constant is 1;
    attribute mti_svvh_generic_type of register_clock_1 : constant is 1;
    attribute mti_svvh_generic_type of register_aclr_1 : constant is 1;
    attribute mti_svvh_generic_type of register_clock_2 : constant is 1;
    attribute mti_svvh_generic_type of register_aclr_2 : constant is 1;
    attribute mti_svvh_generic_type of register_clock_3 : constant is 1;
    attribute mti_svvh_generic_type of register_aclr_3 : constant is 1;
    attribute mti_svvh_generic_type of number_of_multipliers : constant is 1;
    attribute mti_svvh_generic_type of port_sign : constant is 1;
    attribute mti_svvh_generic_type of width_data_in_msb : constant is 3;
    attribute mti_svvh_generic_type of width_data_in_total_msb : constant is 3;
    attribute mti_svvh_generic_type of width_data_out_msb : constant is 3;
    attribute mti_svvh_generic_type of width_data_in_0_msb : constant is 3;
    attribute mti_svvh_generic_type of width_data_in_0_lsb : constant is 1;
    attribute mti_svvh_generic_type of width_data_in_1_msb : constant is 3;
    attribute mti_svvh_generic_type of width_data_in_1_lsb : constant is 3;
    attribute mti_svvh_generic_type of width_data_in_2_msb : constant is 3;
    attribute mti_svvh_generic_type of width_data_in_2_lsb : constant is 3;
    attribute mti_svvh_generic_type of width_data_in_3_msb : constant is 3;
    attribute mti_svvh_generic_type of width_data_in_3_lsb : constant is 3;
end ama_data_split_reg_ext_function;
