library verilog;
use verilog.vl_types.all;
entity common_28nm_ram_block is
    generic(
        operation_mode  : string  := "single_port";
        mixed_port_feed_through_mode: string  := "dont_care";
        init_file_layout: string  := "none";
        ecc_pipeline_stage_enabled: string  := "false";
        enable_ecc      : string  := "false";
        width_eccstatus : integer := 2;
        port_a_first_address: integer := 0;
        port_a_last_address: integer := 0;
        port_a_data_out_clear: string  := "none";
        port_a_data_out_clock: string  := "none";
        port_a_data_width: integer := 1;
        port_a_address_width: integer := 1;
        port_a_byte_enable_mask_width: integer := 1;
        port_b_first_address: integer := 0;
        port_b_last_address: integer := 0;
        port_b_address_clear: string  := "none";
        port_b_data_out_clear: string  := "none";
        port_b_data_in_clock: string  := "clock1";
        port_b_address_clock: string  := "clock1";
        port_b_write_enable_clock: string  := "clock1";
        port_b_read_enable_clock: string  := "clock1";
        port_b_byte_enable_clock: string  := "clock1";
        port_b_data_out_clock: string  := "none";
        port_b_data_width: integer := 1;
        port_b_address_width: integer := 1;
        port_b_byte_enable_mask_width: integer := 1;
        power_up_uninitialized: string  := "false";
        mem_init0       : string  := "";
        mem_init1       : string  := "";
        mem_init2       : string  := "";
        mem_init3       : string  := "";
        mem_init4       : string  := "";
        mem_init5       : string  := "";
        mem_init6       : string  := "";
        mem_init7       : string  := "";
        mem_init8       : string  := "";
        mem_init9       : string  := "";
        clk0_input_clock_enable: string  := "none";
        clk0_core_clock_enable: string  := "none";
        clk0_output_clock_enable: string  := "none";
        clk1_input_clock_enable: string  := "none";
        clk1_core_clock_enable: string  := "none";
        clk1_output_clock_enable: string  := "none";
        bist_ena        : string  := "false";
        port_a_address_clear: string  := "none";
        port_a_write_enable_clock: string  := "clock0";
        port_a_read_enable_clock: string  := "clock0";
        primary_port_is_a: vl_notype;
        primary_port_is_b: vl_notype;
        mode_is_dp      : vl_notype;
        mode_is_sp      : vl_notype;
        mode_is_rom     : vl_notype;
        mode_is_bdp     : vl_notype;
        mode_is_rom_or_sp: vl_notype;
        mixed_port_rdw_is_dont_care: vl_notype;
        out_a_is_reg    : vl_notype;
        out_b_is_reg    : vl_notype;
        data_width      : vl_notype;
        data_unit_width : vl_notype;
        address_width   : vl_notype;
        address_unit_width: vl_notype;
        wired_mode      : vl_notype;
        num_rows        : vl_notype;
        num_cols        : vl_notype;
        mask_width_prime: vl_notype;
        mask_width_sec  : vl_notype;
        byte_size_a     : vl_notype;
        byte_size_b     : vl_notype;
        dual_clock      : vl_notype;
        hw_write_mode_a : vl_notype;
        hw_write_mode_b : vl_notype;
        delay_write_pulse_a: vl_notype;
        delay_write_pulse_b: vl_notype
    );
    port(
        portadatain     : in     vl_logic_vector;
        portaaddr       : in     vl_logic_vector;
        portawe         : in     vl_logic;
        portare         : in     vl_logic;
        portbdatain     : in     vl_logic_vector;
        portbaddr       : in     vl_logic_vector;
        portbwe         : in     vl_logic;
        portbre         : in     vl_logic;
        clk0            : in     vl_logic;
        clk1            : in     vl_logic;
        ena0            : in     vl_logic;
        ena1            : in     vl_logic;
        ena2            : in     vl_logic;
        ena3            : in     vl_logic;
        clr0            : in     vl_logic;
        clr1            : in     vl_logic;
        nerror          : in     vl_logic;
        portabyteenamasks: in     vl_logic_vector;
        portbbyteenamasks: in     vl_logic_vector;
        portaaddrstall  : in     vl_logic;
        portbaddrstall  : in     vl_logic;
        devclrn         : in     vl_logic;
        devpor          : in     vl_logic;
        eccstatus       : out    vl_logic_vector;
        portadataout    : out    vl_logic_vector;
        portbdataout    : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of operation_mode : constant is 1;
    attribute mti_svvh_generic_type of mixed_port_feed_through_mode : constant is 1;
    attribute mti_svvh_generic_type of init_file_layout : constant is 1;
    attribute mti_svvh_generic_type of ecc_pipeline_stage_enabled : constant is 1;
    attribute mti_svvh_generic_type of enable_ecc : constant is 1;
    attribute mti_svvh_generic_type of width_eccstatus : constant is 1;
    attribute mti_svvh_generic_type of port_a_first_address : constant is 1;
    attribute mti_svvh_generic_type of port_a_last_address : constant is 1;
    attribute mti_svvh_generic_type of port_a_data_out_clear : constant is 1;
    attribute mti_svvh_generic_type of port_a_data_out_clock : constant is 1;
    attribute mti_svvh_generic_type of port_a_data_width : constant is 1;
    attribute mti_svvh_generic_type of port_a_address_width : constant is 1;
    attribute mti_svvh_generic_type of port_a_byte_enable_mask_width : constant is 1;
    attribute mti_svvh_generic_type of port_b_first_address : constant is 1;
    attribute mti_svvh_generic_type of port_b_last_address : constant is 1;
    attribute mti_svvh_generic_type of port_b_address_clear : constant is 1;
    attribute mti_svvh_generic_type of port_b_data_out_clear : constant is 1;
    attribute mti_svvh_generic_type of port_b_data_in_clock : constant is 1;
    attribute mti_svvh_generic_type of port_b_address_clock : constant is 1;
    attribute mti_svvh_generic_type of port_b_write_enable_clock : constant is 1;
    attribute mti_svvh_generic_type of port_b_read_enable_clock : constant is 1;
    attribute mti_svvh_generic_type of port_b_byte_enable_clock : constant is 1;
    attribute mti_svvh_generic_type of port_b_data_out_clock : constant is 1;
    attribute mti_svvh_generic_type of port_b_data_width : constant is 1;
    attribute mti_svvh_generic_type of port_b_address_width : constant is 1;
    attribute mti_svvh_generic_type of port_b_byte_enable_mask_width : constant is 1;
    attribute mti_svvh_generic_type of power_up_uninitialized : constant is 1;
    attribute mti_svvh_generic_type of mem_init0 : constant is 1;
    attribute mti_svvh_generic_type of mem_init1 : constant is 1;
    attribute mti_svvh_generic_type of mem_init2 : constant is 1;
    attribute mti_svvh_generic_type of mem_init3 : constant is 1;
    attribute mti_svvh_generic_type of mem_init4 : constant is 1;
    attribute mti_svvh_generic_type of mem_init5 : constant is 1;
    attribute mti_svvh_generic_type of mem_init6 : constant is 1;
    attribute mti_svvh_generic_type of mem_init7 : constant is 1;
    attribute mti_svvh_generic_type of mem_init8 : constant is 1;
    attribute mti_svvh_generic_type of mem_init9 : constant is 1;
    attribute mti_svvh_generic_type of clk0_input_clock_enable : constant is 1;
    attribute mti_svvh_generic_type of clk0_core_clock_enable : constant is 1;
    attribute mti_svvh_generic_type of clk0_output_clock_enable : constant is 1;
    attribute mti_svvh_generic_type of clk1_input_clock_enable : constant is 1;
    attribute mti_svvh_generic_type of clk1_core_clock_enable : constant is 1;
    attribute mti_svvh_generic_type of clk1_output_clock_enable : constant is 1;
    attribute mti_svvh_generic_type of bist_ena : constant is 1;
    attribute mti_svvh_generic_type of port_a_address_clear : constant is 1;
    attribute mti_svvh_generic_type of port_a_write_enable_clock : constant is 1;
    attribute mti_svvh_generic_type of port_a_read_enable_clock : constant is 1;
    attribute mti_svvh_generic_type of primary_port_is_a : constant is 3;
    attribute mti_svvh_generic_type of primary_port_is_b : constant is 3;
    attribute mti_svvh_generic_type of mode_is_dp : constant is 3;
    attribute mti_svvh_generic_type of mode_is_sp : constant is 3;
    attribute mti_svvh_generic_type of mode_is_rom : constant is 3;
    attribute mti_svvh_generic_type of mode_is_bdp : constant is 3;
    attribute mti_svvh_generic_type of mode_is_rom_or_sp : constant is 3;
    attribute mti_svvh_generic_type of mixed_port_rdw_is_dont_care : constant is 3;
    attribute mti_svvh_generic_type of out_a_is_reg : constant is 3;
    attribute mti_svvh_generic_type of out_b_is_reg : constant is 3;
    attribute mti_svvh_generic_type of data_width : constant is 3;
    attribute mti_svvh_generic_type of data_unit_width : constant is 3;
    attribute mti_svvh_generic_type of address_width : constant is 3;
    attribute mti_svvh_generic_type of address_unit_width : constant is 3;
    attribute mti_svvh_generic_type of wired_mode : constant is 3;
    attribute mti_svvh_generic_type of num_rows : constant is 3;
    attribute mti_svvh_generic_type of num_cols : constant is 3;
    attribute mti_svvh_generic_type of mask_width_prime : constant is 3;
    attribute mti_svvh_generic_type of mask_width_sec : constant is 3;
    attribute mti_svvh_generic_type of byte_size_a : constant is 3;
    attribute mti_svvh_generic_type of byte_size_b : constant is 3;
    attribute mti_svvh_generic_type of dual_clock : constant is 3;
    attribute mti_svvh_generic_type of hw_write_mode_a : constant is 3;
    attribute mti_svvh_generic_type of hw_write_mode_b : constant is 3;
    attribute mti_svvh_generic_type of delay_write_pulse_a : constant is 3;
    attribute mti_svvh_generic_type of delay_write_pulse_b : constant is 3;
end common_28nm_ram_block;
