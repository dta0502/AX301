library verilog;
use verilog.vl_types.all;
entity lut_output is
    port(
        \in\            : in     vl_logic;
        \out\           : out    vl_logic
    );
end lut_output;
