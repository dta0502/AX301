library verilog;
use verilog.vl_types.all;
entity cycloneive_routing_wire is
    port(
        datain          : in     vl_logic;
        dataout         : out    vl_logic
    );
end cycloneive_routing_wire;
