library verilog;
use verilog.vl_types.all;
entity row_global is
    port(
        \in\            : in     vl_logic;
        \out\           : out    vl_logic
    );
end row_global;
