library verilog;
use verilog.vl_types.all;
entity PRIM_GDFF_LOW is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end PRIM_GDFF_LOW;
