library verilog;
use verilog.vl_types.all;
entity opndrn is
    port(
        \in\            : in     vl_logic;
        \out\           : out    vl_logic
    );
end opndrn;
